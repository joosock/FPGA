module ex_multiplier(a,b,m);

input [3:0] a;
input [3:0] b;

output [7:0] m;

assign m = a*b; 

endmodule